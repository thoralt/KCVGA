LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SyncGenerator IS GENERIC
(
    H_TOTAL, V_TOTAL, V_ACTIVE_END, H_SYNC_PULSE_LENGTH, V_SYNC_PULSE_LENGTH : NATURAL;
    H_POLARITY, V_POLARITY                                                   : STD_LOGIC
);
PORT
(
    HPOS      : INTEGER RANGE 0 TO H_TOTAL - 1;
    VPOS      : INTEGER RANGE 0 TO V_TOTAL - 1;
    HSYNC     : OUT STD_LOGIC;
    VSYNC     : OUT STD_LOGIC;
    FRAMESYNC : OUT STD_LOGIC
);
END SyncGenerator;

ARCHITECTURE Behavioral OF SyncGenerator IS

BEGIN

    HSYNC <= H_POLARITY WHEN HPOS < H_SYNC_PULSE_LENGTH ELSE
        NOT H_POLARITY;
    VSYNC <= V_POLARITY WHEN VPOS < V_SYNC_PULSE_LENGTH ELSE
        NOT V_POLARITY;
    FRAMESYNC <= '1' WHEN VPOS = V_ACTIVE_END ELSE
        '0';

END Behavioral;
